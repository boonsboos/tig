module main

fn main() {
	println('hello world')

	// autosave thread
	// game thread	
}