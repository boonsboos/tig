module graphics

import term.ui

pub fn draw_money_rectangle() {

}