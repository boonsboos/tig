module main

import util

__global options = util.parse_args()

fn main() {
	println(options)
	// autosave thread
	// game thread	
}