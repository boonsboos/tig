module game

import term

fn handle_input() {
	
}