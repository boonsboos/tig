module main

fn main()
{
	println('hello world')	
}